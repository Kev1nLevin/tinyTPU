/home/kevinlevin/Projects/Neural_Network_Accelerator/techlef/asap7_tech_4x_201209.lef