// =============================================================================
// Module: activation_unit
// Description: Configurable activation function unit (Production)
//              Replaces gelu_unit with multi-function support.
//
//              Supported functions (selected by act_func):
//                3'b000 = NONE  (passthrough)
//                3'b001 = ReLU  (max(0, x))
//                3'b010 = GeLU  (256-entry hardcoded LUT, x ∈ [-4, +4))
//
//              Hardcoded 256-entry FP32 LUT (no $readmemh — synthesis clean).
//              x ≤ -4 → 0.0  |  x ≥ +4 → x (passthrough)
//
//              Output is REGISTERED for timing closure.
// =============================================================================

module activation_unit (
    input  logic        clk,
    input  logic        rst_n,
    input  logic        valid_in,   // pulse: data is valid, capture output
    input  logic [31:0] fp32_in,    // FP32 input value
    input  logic [2:0]  act_func,   // activation function select
    input  logic [31:0] bias_val,   // FP32 bias to add (0 if disabled)
    input  logic        bias_en,    // 1 = add bias before activation
    output logic [31:0] fp32_out,   // FP32 result (registered)
    output logic        valid_out   // delayed valid
);

    // =========================================================================
    // Activation function encoding
    // =========================================================================
    localparam [2:0] ACT_NONE = 3'b000;
    localparam [2:0] ACT_RELU = 3'b001;
    localparam [2:0] ACT_GELU = 3'b010;

    // =========================================================================
    // FP32 field extraction (from input, used for LUT addressing and ReLU)
    // =========================================================================
    logic        fp_sign;
    logic [7:0]  fp_exp;
    logic [22:0] fp_mant;

    assign fp_sign = fp32_in[31];
    assign fp_exp  = fp32_in[30:23];
    assign fp_mant = fp32_in[22:0];

    // |x| >= 4.0 check (biased exp >= 129)
    logic abs_ge_4;
    assign abs_ge_4 = (fp_exp >= 8'd129);

    // =========================================================================
    // GeLU LUT address computation (same as original gelu_unit)
    // =========================================================================
    logic [6:0] mag_idx;

    always_comb begin
        case (fp_exp)
            8'd128:  mag_idx = {1'b1,    fp_mant[22:17]};
            8'd127:  mag_idx = {2'b01,   fp_mant[22:18]};
            8'd126:  mag_idx = {3'b001,  fp_mant[22:19]};
            8'd125:  mag_idx = {4'b0001, fp_mant[22:20]};
            8'd124:  mag_idx = {5'b00001,fp_mant[22:21]};
            8'd123:  mag_idx = {6'b000001,fp_mant[22]};
            default: mag_idx = 7'd0;
        endcase
    end

    logic [7:0] lut_addr;
    always_comb begin
        if (abs_ge_4)     lut_addr = 8'd0;
        else if (fp_sign) lut_addr = 8'd128 - {1'b0, mag_idx};
        else              lut_addr = 8'd128 + {1'b0, mag_idx};
    end

    // =========================================================================
    // Hardcoded 256-entry GeLU LUT (synthesis-clean, no $readmemh)
    // Generated by: x = (i-128)/32; GeLU(x) = x*0.5*(1+tanh(0.7978846*(x+0.044715*x³)))
    // =========================================================================
    logic [31:0] lut_data;

    always_comb begin
        case (lut_addr)
            8'd0: lut_data = 32'hB89350FC;
            8'd1: lut_data = 32'hB8AADA4F;
            8'd2: lut_data = 32'hB8C5CF05;
            8'd3: lut_data = 32'hB8E4A052;
            8'd4: lut_data = 32'hB903E5FE;
            8'd5: lut_data = 32'hB917EEBB;
            8'd6: lut_data = 32'hB92EB78C;
            8'd7: lut_data = 32'hB94895A9;
            8'd8: lut_data = 32'hB965E700;
            8'd9: lut_data = 32'hB9838973;
            8'd10: lut_data = 32'hB9964567;
            8'd11: lut_data = 32'hB9AB657F;
            8'd12: lut_data = 32'hB9C32DB3;
            8'd13: lut_data = 32'hB9DDE82B;
            8'd14: lut_data = 32'hB9FBE5B2;
            8'd15: lut_data = 32'hBA0EBF0B;
            8'd16: lut_data = 32'hBA21884F;
            8'd17: lut_data = 32'hBA368237;
            8'd18: lut_data = 32'hBA4DE480;
            8'd19: lut_data = 32'hBA67EB44;
            8'd20: lut_data = 32'hBA826B9A;
            8'd21: lut_data = 32'hBA9276E8;
            8'd22: lut_data = 32'hBAA43CC9;
            8'd23: lut_data = 32'hBAB7E518;
            8'd24: lut_data = 32'hBACD9A60;
            8'd25: lut_data = 32'hBAE589F4;
            8'd26: lut_data = 32'hBAFFE408;
            8'd27: lut_data = 32'hBB0E6DE1;
            8'd28: lut_data = 32'hBB1E53A4;
            8'd29: lut_data = 32'hBB2FBFEA;
            8'd30: lut_data = 32'hBB42D0DC;
            8'd31: lut_data = 32'hBB57A637;
            8'd32: lut_data = 32'hBB6E614B;
            8'd33: lut_data = 32'hBB83927E;
            8'd34: lut_data = 32'hBB910ADF;
            8'd35: lut_data = 32'hBB9FACCA;
            8'd36: lut_data = 32'hBBAF8C02;
            8'd37: lut_data = 32'hBBC0BD07;
            8'd38: lut_data = 32'hBBD35511;
            8'd39: lut_data = 32'hBBE76A04;
            8'd40: lut_data = 32'hBBFD1269;
            8'd41: lut_data = 32'hBC0A32B0;
            8'd42: lut_data = 32'hBC16BD49;
            8'd43: lut_data = 32'hBC243511;
            8'd44: lut_data = 32'hBC32A64F;
            8'd45: lut_data = 32'hBC421D70;
            8'd46: lut_data = 32'hBC52A703;
            8'd47: lut_data = 32'hBC644FA6;
            8'd48: lut_data = 32'hBC7723FB;
            8'd49: lut_data = 32'hBC85984E;
            8'd50: lut_data = 32'hBC904102;
            8'd51: lut_data = 32'hBC9B9242;
            8'd52: lut_data = 32'hBCA79217;
            8'd53: lut_data = 32'hBCB4465F;
            8'd54: lut_data = 32'hBCC1B4C5;
            8'd55: lut_data = 32'hBCCFE2B6;
            8'd56: lut_data = 32'hBCDED550;
            8'd57: lut_data = 32'hBCEE915C;
            8'd58: lut_data = 32'hBCFF1B3E;
            8'd59: lut_data = 32'hBD083B73;
            8'd60: lut_data = 32'hBD1153E4;
            8'd61: lut_data = 32'hBD1AD861;
            8'd62: lut_data = 32'hBD24CA0D;
            8'd63: lut_data = 32'hBD2F29B4;
            8'd64: lut_data = 32'hBD39F7C2;
            8'd65: lut_data = 32'hBD45343E;
            8'd66: lut_data = 32'hBD50DEBF;
            8'd67: lut_data = 32'hBD5CF666;
            8'd68: lut_data = 32'hBD6979D5;
            8'd69: lut_data = 32'hBD766727;
            8'd70: lut_data = 32'hBD81DDF3;
            8'd71: lut_data = 32'hBD88BA83;
            8'd72: lut_data = 32'hBD8FC76F;
            8'd73: lut_data = 32'hBD97028C;
            8'd74: lut_data = 32'hBD9E695B;
            8'd75: lut_data = 32'hBDA5F8FF;
            8'd76: lut_data = 32'hBDADAE41;
            8'd77: lut_data = 32'hBDB58585;
            8'd78: lut_data = 32'hBDBD7ACC;
            8'd79: lut_data = 32'hBDC589B3;
            8'd80: lut_data = 32'hBDCDAD69;
            8'd81: lut_data = 32'hBDD5E0B7;
            8'd82: lut_data = 32'hBDDE1DF6;
            8'd83: lut_data = 32'hBDE65F13;
            8'd84: lut_data = 32'hBDEE9D8C;
            8'd85: lut_data = 32'hBDF6D272;
            8'd86: lut_data = 32'hBDFEF665;
            8'd87: lut_data = 32'hBE0380CD;
            8'd88: lut_data = 32'hBE0775ED;
            8'd89: lut_data = 32'hBE0B5640;
            8'd90: lut_data = 32'hBE0F1D40;
            8'd91: lut_data = 32'hBE12C638;
            8'd92: lut_data = 32'hBE164C3D;
            8'd93: lut_data = 32'hBE19AA39;
            8'd94: lut_data = 32'hBE1CDAEA;
            8'd95: lut_data = 32'hBE1FD8E2;
            8'd96: lut_data = 32'hBE229E90;
            8'd97: lut_data = 32'hBE25263E;
            8'd98: lut_data = 32'hBE276A17;
            8'd99: lut_data = 32'hBE29642C;
            8'd100: lut_data = 32'hBE2B0E73;
            8'd101: lut_data = 32'hBE2C62D4;
            8'd102: lut_data = 32'hBE2D5B26;
            8'd103: lut_data = 32'hBE2DF137;
            8'd104: lut_data = 32'hBE2E1ED1;
            8'd105: lut_data = 32'hBE2DDDC1;
            8'd106: lut_data = 32'hBE2D27D7;
            8'd107: lut_data = 32'hBE2BF6F2;
            8'd108: lut_data = 32'hBE2A4500;
            8'd109: lut_data = 32'hBE280C0A;
            8'd110: lut_data = 32'hBE254633;
            8'd111: lut_data = 32'hBE21EDC2;
            8'd112: lut_data = 32'hBE1DFD25;
            8'd113: lut_data = 32'hBE196EFB;
            8'd114: lut_data = 32'hBE143E15;
            8'd115: lut_data = 32'hBE0E657C;
            8'd116: lut_data = 32'hBE07E079;
            8'd117: lut_data = 32'hBE00AA97;
            8'd118: lut_data = 32'hBDF17F54;
            8'd119: lut_data = 32'hBDE037A5;
            8'd120: lut_data = 32'hBDCD7702;
            8'd121: lut_data = 32'hBDB936F8;
            8'd122: lut_data = 32'hBDA371C3;
            8'd123: lut_data = 32'hBD8C2258;
            8'd124: lut_data = 32'hBD6688CB;
            8'd125: lut_data = 32'hBD31A8C1;
            8'd126: lut_data = 32'hBCF33E00;
            8'd127: lut_data = 32'hBC799E33;
            8'd128: lut_data = 32'h00000000;
            8'd129: lut_data = 32'h3C8330E6;
            8'd130: lut_data = 32'h3D066100;
            8'd131: lut_data = 32'h3D4E573F;
            8'd132: lut_data = 32'h3D8CBB9A;
            8'd133: lut_data = 32'h3DB3DDA8;
            8'd134: lut_data = 32'h3DDC8E3D;
            8'd135: lut_data = 32'h3E036484;
            8'd136: lut_data = 32'h3E19447F;
            8'd137: lut_data = 32'h3E2FE42E;
            8'd138: lut_data = 32'h3E474056;
            8'd139: lut_data = 32'h3E5F5569;
            8'd140: lut_data = 32'h3E781F87;
            8'd141: lut_data = 32'h3E88CD42;
            8'd142: lut_data = 32'h3E95E0F6;
            8'd143: lut_data = 32'h3EA34882;
            8'd144: lut_data = 32'h3EB1016D;
            8'd145: lut_data = 32'h3EBF091F;
            8'd146: lut_data = 32'h3ECD5CE7;
            8'd147: lut_data = 32'h3EDBF9FB;
            8'd148: lut_data = 32'h3EEADD80;
            8'd149: lut_data = 32'h3EFA0487;
            8'd150: lut_data = 32'h3F04B60A;
            8'd151: lut_data = 32'h3F0C8890;
            8'd152: lut_data = 32'h3F14784C;
            8'd153: lut_data = 32'h3F1C83B2;
            8'd154: lut_data = 32'h3F24A937;
            8'd155: lut_data = 32'h3F2CE74B;
            8'd156: lut_data = 32'h3F353C63;
            8'd157: lut_data = 32'h3F3DA6F5;
            8'd158: lut_data = 32'h3F46257A;
            8'd159: lut_data = 32'h3F4EB670;
            8'd160: lut_data = 32'h3F57585C;
            8'd161: lut_data = 32'h3F6009C7;
            8'd162: lut_data = 32'h3F68C946;
            8'd163: lut_data = 32'h3F719572;
            8'd164: lut_data = 32'h3F7A6CF1;
            8'd165: lut_data = 32'h3F81A739;
            8'd166: lut_data = 32'h3F861C58;
            8'd167: lut_data = 32'h3F8A9538;
            8'd168: lut_data = 32'h3F8F1142;
            8'd169: lut_data = 32'h3F938FE6;
            8'd170: lut_data = 32'h3F98109A;
            8'd171: lut_data = 32'h3F9C92D9;
            8'd172: lut_data = 32'h3FA11627;
            8'd173: lut_data = 32'h3FA59A0F;
            8'd174: lut_data = 32'h3FAA1E21;
            8'd175: lut_data = 32'h3FAEA1F5;
            8'd176: lut_data = 32'h3FB32529;
            8'd177: lut_data = 32'h3FB7A765;
            8'd178: lut_data = 32'h3FBC2853;
            8'd179: lut_data = 32'h3FC0A7A8;
            8'd180: lut_data = 32'h3FC5251C;
            8'd181: lut_data = 32'h3FC9A070;
            8'd182: lut_data = 32'h3FCE196A;
            8'd183: lut_data = 32'h3FD28FD7;
            8'd184: lut_data = 32'h3FD70389;
            8'd185: lut_data = 32'h3FDB7458;
            8'd186: lut_data = 32'h3FDFE221;
            8'd187: lut_data = 32'h3FE44CC7;
            8'd188: lut_data = 32'h3FE8B431;
            8'd189: lut_data = 32'h3FED184D;
            8'd190: lut_data = 32'h3FF1790A;
            8'd191: lut_data = 32'h3FF5D65E;
            8'd192: lut_data = 32'h3FFA3042;
            8'd193: lut_data = 32'h3FFE86B2;
            8'd194: lut_data = 32'h40016CD8;
            8'd195: lut_data = 32'h4003949E;
            8'd196: lut_data = 32'h4005BAB0;
            8'd197: lut_data = 32'h4007DF12;
            8'd198: lut_data = 32'h400A01CA;
            8'd199: lut_data = 32'h400C22DD;
            8'd200: lut_data = 32'h400E4255;
            8'd201: lut_data = 32'h4010603B;
            8'd202: lut_data = 32'h40127C96;
            8'd203: lut_data = 32'h40149773;
            8'd204: lut_data = 32'h4016B0DC;
            8'd205: lut_data = 32'h4018C8DB;
            8'd206: lut_data = 32'h401ADF7E;
            8'd207: lut_data = 32'h401CF4CF;
            8'd208: lut_data = 32'h401F08DC;
            8'd209: lut_data = 32'h40211BB0;
            8'd210: lut_data = 32'h40232D59;
            8'd211: lut_data = 32'h40253DE3;
            8'd212: lut_data = 32'h40274D5A;
            8'd213: lut_data = 32'h40295BCB;
            8'd214: lut_data = 32'h402B6943;
            8'd215: lut_data = 32'h402D75CD;
            8'd216: lut_data = 32'h402F8177;
            8'd217: lut_data = 32'h40318C4B;
            8'd218: lut_data = 32'h40339655;
            8'd219: lut_data = 32'h40359FA1;
            8'd220: lut_data = 32'h4037A83A;
            8'd221: lut_data = 32'h4039B02A;
            8'd222: lut_data = 32'h403BB77B;
            8'd223: lut_data = 32'h403DBE37;
            8'd224: lut_data = 32'h403FC468;
            8'd225: lut_data = 32'h4041CA16;
            8'd226: lut_data = 32'h4043CF4C;
            8'd227: lut_data = 32'h4045D410;
            8'd228: lut_data = 32'h4047D86B;
            8'd229: lut_data = 32'h4049DC65;
            8'd230: lut_data = 32'h404BE003;
            8'd231: lut_data = 32'h404DE34F;
            8'd232: lut_data = 32'h404FE64D;
            8'd233: lut_data = 32'h4051E903;
            8'd234: lut_data = 32'h4053EB78;
            8'd235: lut_data = 32'h4055EDB1;
            8'd236: lut_data = 32'h4057EFB3;
            8'd237: lut_data = 32'h4059F181;
            8'd238: lut_data = 32'h405BF322;
            8'd239: lut_data = 32'h405DF498;
            8'd240: lut_data = 32'h405FF5E7;
            8'd241: lut_data = 32'h4061F714;
            8'd242: lut_data = 32'h4063F821;
            8'd243: lut_data = 32'h4065F911;
            8'd244: lut_data = 32'h4067F9E7;
            8'd245: lut_data = 32'h4069FAA5;
            8'd246: lut_data = 32'h406BFB4E;
            8'd247: lut_data = 32'h406DFBE4;
            8'd248: lut_data = 32'h406FFC68;
            8'd249: lut_data = 32'h4071FCDE;
            8'd250: lut_data = 32'h4073FD45;
            8'd251: lut_data = 32'h4075FDA0;
            8'd252: lut_data = 32'h4077FDF0;
            8'd253: lut_data = 32'h4079FE37;
            8'd254: lut_data = 32'h407BFE74;
            8'd255: lut_data = 32'h407DFEAA;
            default: lut_data = 32'h00000000;
        endcase
    end

    // =========================================================================
    // Activation function MUX (combinational)
    // =========================================================================
    logic [31:0] act_result;

    always_comb begin
        case (act_func)
            ACT_NONE: begin
                act_result = fp32_in;
            end

            ACT_RELU: begin
                // ReLU: max(0, x) — just check sign bit
                act_result = fp_sign ? 32'h0000_0000 : fp32_in;
            end

            ACT_GELU: begin
                if (abs_ge_4 && fp_sign)
                    act_result = 32'h0000_0000;     // x <= -4 → 0
                else if (abs_ge_4 && !fp_sign)
                    act_result = fp32_in;            // x >= +4 → x
                else
                    act_result = lut_data;
            end

            default: begin
                act_result = fp32_in;  // unknown → passthrough
            end
        endcase
    end

    // =========================================================================
    // Output register (breaks timing-critical path)
    // =========================================================================
    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            fp32_out  <= '0;
            valid_out <= 1'b0;
        end else begin
            valid_out <= valid_in;
            if (valid_in)
                fp32_out <= act_result;
        end
    end

endmodule
