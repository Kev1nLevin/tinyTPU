/home/kevinlevin/Projects/Neural_Network_Accelerator/lef/scaled/asap7sc7p5t_28_L_4x_220121a.lef